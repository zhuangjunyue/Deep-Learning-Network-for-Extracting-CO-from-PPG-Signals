module LAYER3(
    input clk,
    input reset,
    input valid_in, // 上游模块数据有效信号
    input logic signed[15:0] input_data[0:31], // 32个Q4.12格式的输入数据
    output logic signed[15:0] output_data[0:15], // 16个Q4.12格式的输出数据
    output logic valid_out, // 输出数据有效信号
    output ready_out // 准备好接收下游数据的信号
);


// 定义一个16位宽有符号整数的32元素一维数组类型
typedef logic signed [15:0] signed_matrix_1x32_t[32];

// 定义一个此类型的16元素一维数组，即16x32的二维数组
typedef signed_matrix_1x32_t signed_matrix_16x32_t[16];


const signed_matrix_16x32_t weights_3 = '{

'{-16'sd652, -16'sd1112, -16'sd413, -16'sd118, 16'sd1429, 16'sd1181, -16'sd1028, 16'sd381, 16'sd370, 16'sd654, 16'sd174, 16'sd1912, -16'sd322, 16'sd736, 16'sd1194, 16'sd126, -16'sd566, -16'sd1393, 16'sd1404, -16'sd504, -16'sd105, 16'sd243, -16'sd1201, 16'sd828, -16'sd629, 16'sd64, -16'sd446, -16'sd439, 16'sd323, -16'sd752, -16'sd1299, 16'sd754},
'{16'sd334, -16'sd252, -16'sd764, 16'sd636, -16'sd1390, 16'sd775, 16'sd2801, -16'sd969, -16'sd1475, 16'sd190, -16'sd597, -16'sd40, -16'sd39, 16'sd1202, -16'sd1235, -16'sd1054, -16'sd1514, -16'sd397, -16'sd646, 16'sd2220, -16'sd648, 16'sd214, 16'sd97, 16'sd732, -16'sd547, 16'sd2054, -16'sd59, -16'sd2067, 16'sd753, -16'sd1044, 16'sd453, 16'sd1688},
'{16'sd1161, 16'sd18, -16'sd801, 16'sd90, 16'sd1535, 16'sd1793, 16'sd202, 16'sd355, -16'sd122, -16'sd591, 16'sd989, 16'sd182, 16'sd189, -16'sd618, 16'sd887, 16'sd599, -16'sd26, -16'sd294, -16'sd1229, -16'sd101, -16'sd247, -16'sd688, -16'sd638, -16'sd500, -16'sd1760, -16'sd2090, 16'sd263, 16'sd1147, -16'sd210, 16'sd1173, -16'sd315, 16'sd126},
'{16'sd1943, -16'sd1421, 16'sd522, 16'sd382, 16'sd768, 16'sd382, 16'sd636, 16'sd1850, -16'sd1280, 16'sd724, -16'sd629, 16'sd107, 16'sd486, 16'sd646, -16'sd718, -16'sd207, -16'sd243, 16'sd904, 16'sd1372, -16'sd1868, 16'sd750, 16'sd715, -16'sd60, -16'sd1913, -16'sd1975, -16'sd1769, -16'sd136, -16'sd173, 16'sd1312, -16'sd837, 16'sd295, -16'sd613},
'{-16'sd381, -16'sd700, -16'sd1088, 16'sd1042, 16'sd761, 16'sd803, -16'sd1862, 16'sd531, 16'sd395, 16'sd1173, 16'sd395, 16'sd1188, 16'sd1339, 16'sd1900, 16'sd789, -16'sd642, 16'sd759, -16'sd649, 16'sd796, 16'sd356, -16'sd382, -16'sd1226, -16'sd716, 16'sd108, -16'sd402, -16'sd1038, -16'sd2251, 16'sd1397, 16'sd500, 16'sd5, -16'sd571, -16'sd241},
'{-16'sd1122, -16'sd418, 16'sd770, -16'sd313, -16'sd704, -16'sd197, 16'sd158, -16'sd1085, -16'sd924, 16'sd746, 16'sd1343, -16'sd2413, 16'sd54, 16'sd583, -16'sd66, -16'sd611, 16'sd3556, 16'sd742, 16'sd916, -16'sd862, 16'sd232, 16'sd46, 16'sd1024, 16'sd2729, 16'sd856, -16'sd425, -16'sd517, -16'sd104, 16'sd884, -16'sd2012, -16'sd448, 16'sd737},
'{16'sd765, -16'sd758, -16'sd1313, -16'sd1748, -16'sd552, 16'sd160, -16'sd230, -16'sd455, -16'sd1558, -16'sd1512, 16'sd55, -16'sd296, -16'sd2, 16'sd464, -16'sd1613, -16'sd1054, 16'sd829, -16'sd324, 16'sd488, -16'sd522, -16'sd107, -16'sd312, 16'sd232, 16'sd443, 16'sd1690, -16'sd192, -16'sd415, 16'sd1577, 16'sd411, 16'sd310, -16'sd1193, 16'sd551},
'{16'sd701, -16'sd206, -16'sd237, 16'sd1684, -16'sd149, -16'sd44, 16'sd1295, -16'sd396, -16'sd510, 16'sd646, 16'sd830, 16'sd678, 16'sd786, -16'sd1512, 16'sd55, -16'sd556, 16'sd524, 16'sd1540, -16'sd273, -16'sd670, 16'sd1076, -16'sd817, -16'sd796, -16'sd1562, 16'sd175, 16'sd489, -16'sd1015, -16'sd87, -16'sd299, 16'sd2346, 16'sd712, 16'sd450},
'{16'sd1061, 16'sd1031, -16'sd3601, 16'sd304, -16'sd293, -16'sd473, 16'sd1868, -16'sd775, -16'sd1535, -16'sd1668, -16'sd1312, 16'sd1294, 16'sd520, 16'sd780, -16'sd1541, -16'sd2347, 16'sd527, -16'sd320, 16'sd1767, 16'sd454, 16'sd36, -16'sd1118, -16'sd1049, 16'sd634, 16'sd734, -16'sd767, -16'sd1825, -16'sd1556, -16'sd967, -16'sd900, 16'sd733, -16'sd692},
'{-16'sd99, -16'sd972, -16'sd337, 16'sd235, -16'sd1729, 16'sd1898, 16'sd142, -16'sd852, -16'sd755, -16'sd150, 16'sd130, 16'sd1097, -16'sd757, 16'sd1093, -16'sd1086, 16'sd799, -16'sd1552, 16'sd1885, -16'sd872, 16'sd987, -16'sd1685, 16'sd1264, 16'sd67, 16'sd1572, -16'sd393, 16'sd1105, 16'sd2592, -16'sd51, 16'sd1383, -16'sd833, -16'sd833, -16'sd180},
'{-16'sd78, -16'sd385, -16'sd278, -16'sd1642, 16'sd75, -16'sd215, 16'sd245, 16'sd803, 16'sd93, -16'sd900, 16'sd2320, -16'sd1507, -16'sd741, -16'sd211, 16'sd1176, -16'sd1156, -16'sd1230, 16'sd489, 16'sd383, 16'sd165, 16'sd1074, 16'sd1138, -16'sd483, -16'sd1733, -16'sd804, -16'sd1645, -16'sd1156, 16'sd1193, 16'sd812, 16'sd986, 16'sd1135, 16'sd1051},
'{16'sd278, -16'sd237, 16'sd1066, 16'sd333, 16'sd913, 16'sd277, 16'sd275, 16'sd399, -16'sd114, 16'sd256, -16'sd143, -16'sd808, -16'sd1565, 16'sd797, 16'sd1690, 16'sd1694, 16'sd763, 16'sd926, 16'sd2460, -16'sd448, 16'sd1286, 16'sd770, -16'sd1145, -16'sd1563, -16'sd820, -16'sd1010, -16'sd362, -16'sd1358, 16'sd46, 16'sd668, -16'sd534, -16'sd847},
'{16'sd1410, -16'sd638, 16'sd2364, 16'sd563, -16'sd63, 16'sd758, -16'sd892, 16'sd710, 16'sd1187, -16'sd1323, 16'sd192, 16'sd1415, 16'sd3263, -16'sd2407, 16'sd2143, -16'sd993, -16'sd1131, 16'sd1261, 16'sd952, -16'sd487, -16'sd341, 16'sd355, 16'sd830, 16'sd1740, -16'sd1350, -16'sd1964, -16'sd1700, -16'sd263, -16'sd1171, -16'sd368, 16'sd330, -16'sd1843},
'{-16'sd916, 16'sd490, -16'sd207, 16'sd1211, -16'sd1046, 16'sd1668, 16'sd280, -16'sd730, 16'sd982, 16'sd1062, -16'sd945, 16'sd147, 16'sd170, -16'sd1266, 16'sd1622, -16'sd1534, -16'sd1264, -16'sd289, 16'sd134, -16'sd2347, 16'sd819, -16'sd685, 16'sd880, -16'sd2149, -16'sd742, -16'sd618, -16'sd490, -16'sd1793, 16'sd1362, -16'sd856, 16'sd879, -16'sd614},
'{-16'sd437, 16'sd318, -16'sd770, 16'sd1818, 16'sd279, -16'sd1177, -16'sd130, 16'sd810, -16'sd1297, 16'sd1633, -16'sd1196, -16'sd1647, -16'sd1348, -16'sd474, 16'sd504, 16'sd1015, -16'sd1212, -16'sd856, 16'sd176, -16'sd208, -16'sd310, -16'sd622, -16'sd135, -16'sd1042, -16'sd408, -16'sd1695, 16'sd23, 16'sd2133, 16'sd900, -16'sd475, -16'sd1287, 16'sd412},
'{16'sd39, -16'sd785, -16'sd1072, -16'sd1103, 16'sd1681, -16'sd1087, -16'sd805, 16'sd397, -16'sd803, 16'sd395, -16'sd1158, 16'sd1796, 16'sd340, -16'sd980, -16'sd577, -16'sd488, -16'sd466, -16'sd1678, -16'sd905, -16'sd1828, 16'sd1745, -16'sd24, 16'sd543, 16'sd17, -16'sd314, 16'sd1642, -16'sd424, 16'sd910, -16'sd587, -16'sd952, -16'sd118, -16'sd330  }



};

typedef logic signed [15:0] signed_matrix_1x16_t[16];



const signed_matrix_1x16_t biases_3 = '{-16'sd6, -16'sd7, -16'sd14, 16'sd3, 16'sd1, -16'sd3, -16'sd7, 16'sd3, 16'sd3, 16'sd3, 16'sd9, 16'sd2, 16'sd3, -16'sd2, -16'sd1, 16'sd4};

integer i, j; 
logic signed [31:0] sum; // 用于累加，扩展位宽以避免溢出


logic signed [15:0] temp_output_data[0:15]; // 临时存储调整后的结果

always @(posedge clk or posedge reset) begin
    if (reset) begin
        for (i = 0; i < 16; i = i + 1) begin
            output_data[i] <= 0; // 清零输出数据
        end
        valid_out <= 0; // 重置时输出数据无效
    end else if (valid_in) begin
        for (i = 0; i < 16; i = i + 1) begin
            sum = 0; // 在开始累加前初始化sum为0
            for (j = 0; j < 32; j = j + 1) begin
                // 执行矩阵乘法和累加
                sum = sum + (input_data[j] * weights_3[i][j]);
            end
            // 所有加权和完成后，整体右移12位来调整格式
            sum = sum >>> 12;
            sum = sum + biases_3[i];
            // 临时存储调整后的结果
            temp_output_data[i] = sum[15:0];
        end
        // 统一更新输出数据
        for (i = 0; i < 16; i = i + 1) begin
            output_data[i] <= temp_output_data[i];
        end
        valid_out <= 1; // 处理完成后，标记输出数据为有效
    end
end


assign ready_out = 1;



endmodule
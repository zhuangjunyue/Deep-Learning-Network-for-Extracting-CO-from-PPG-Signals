module LAYER2(
    input clk,
    input reset,
    input valid_in, // 上游模块数据有效信号
    input logic signed[15:0] input_data[0:63], // 64个Q4.12格式的输入数据
    output logic signed[15:0] output_data[0:31], // 32个Q4.12格式的输出数据
    output logic valid_out, // 输出数据有效信号
    output ready_out // 准备好接收下游数据的信号
);
// 假设权重和偏置已经硬编码

typedef logic signed [15:0] signed_matrix_1x64_t[64];

// 定义一个此类型的64元素一维数组，即二维数组
typedef signed_matrix_1x64_t signed_matrix_32x64_t[32];


const signed_matrix_32x64_t weights_2 = '{
   

  


'{16'sd770, -16'sd518, 16'sd178, -16'sd511, 16'sd1143, -16'sd2108, -16'sd23, -16'sd421, 16'sd927, -16'sd76, 16'sd567, -16'sd744, -16'sd539, -16'sd736, -16'sd558, 16'sd1321,16'sd786, 16'sd525, -16'sd169, 16'sd575, -16'sd684, 16'sd1786, -16'sd108, -16'sd151, 16'sd808, -16'sd297, 16'sd1027, -16'sd461, 16'sd233, -16'sd245, -16'sd368, -16'sd326,16'sd127, 16'sd259, -16'sd429, -16'sd119, -16'sd346, -16'sd230, -16'sd1179, -16'sd1012, 16'sd188, -16'sd241, 16'sd23, -16'sd175, 16'sd514, -16'sd272, 16'sd522, -16'sd229,16'sd222, 16'sd462, -16'sd385, 16'sd1404, 16'sd435, 16'sd935, 16'sd951, -16'sd588, 16'sd485, 16'sd49, 16'sd523, -16'sd437, -16'sd395, -16'sd1480, 16'sd215, -16'sd30},
'{16'sd671, 16'sd282, -16'sd152, -16'sd275, 16'sd1614, 16'sd1024, 16'sd628, 16'sd90, -16'sd954, 16'sd753, -16'sd521, -16'sd640, 16'sd1255, -16'sd557, -16'sd543, 16'sd813,16'sd482, -16'sd103, -16'sd619, -16'sd1299, 16'sd719, -16'sd750, 16'sd327, 16'sd420, -16'sd662, 16'sd60, 16'sd177, 16'sd460, 16'sd124, -16'sd838, 16'sd790, 16'sd896,16'sd1057, 16'sd878, -16'sd108, -16'sd962, -16'sd545, -16'sd1526, 16'sd473, 16'sd708, -16'sd907, 16'sd1211, -16'sd1323, 16'sd21, 16'sd794, 16'sd331, -16'sd918, -16'sd1083,16'sd502, 16'sd103, -16'sd271, 16'sd404, 16'sd69, -16'sd352, -16'sd680, -16'sd19, -16'sd815, -16'sd196, -16'sd980, 16'sd567, -16'sd470, 16'sd672, -16'sd1003, -16'sd203},
'{-16'sd139, -16'sd107, 16'sd1084, -16'sd114, -16'sd11, 16'sd659, -16'sd455, -16'sd213, 16'sd255, -16'sd916, 16'sd1756, 16'sd592, -16'sd1087, 16'sd555, -16'sd279, -16'sd79,16'sd478, -16'sd415, -16'sd154, -16'sd624, 16'sd99, -16'sd740, -16'sd405, -16'sd518, 16'sd6, 16'sd370, 16'sd1170, 16'sd396, -16'sd77, -16'sd326, -16'sd1599, -16'sd929,16'sd636, 16'sd759, 16'sd1076, -16'sd637, 16'sd295, -16'sd1658, 16'sd68, 16'sd375, -16'sd114, -16'sd784, 16'sd1257, 16'sd13, 16'sd1126, 16'sd290, -16'sd730, -16'sd390,16'sd1224, 16'sd1020, 16'sd51, 16'sd721, -16'sd455, -16'sd56, 16'sd511, 16'sd791, -16'sd1451, 16'sd61, 16'sd275, -16'sd906, -16'sd333, -16'sd343, -16'sd703, -16'sd46},
'{-16'sd309, 16'sd1172, -16'sd700, 16'sd533, 16'sd638, -16'sd1137, -16'sd403, -16'sd915, 16'sd175, -16'sd645, 16'sd378, 16'sd586, -16'sd776, -16'sd7, 16'sd721, -16'sd104,16'sd657, -16'sd314, -16'sd204, -16'sd847, -16'sd494, -16'sd351, 16'sd958, 16'sd1263, -16'sd1754, -16'sd255, 16'sd82, -16'sd1586, 16'sd428, 16'sd583, 16'sd74, -16'sd816,16'sd1146, -16'sd828, -16'sd1344, -16'sd12, -16'sd283, -16'sd221, -16'sd884, 16'sd1490, 16'sd424, -16'sd976, -16'sd233, 16'sd89, -16'sd599, -16'sd87, 16'sd30, 16'sd1706,16'sd435, 16'sd45, -16'sd186, 16'sd781, 16'sd761, -16'sd933, -16'sd280, 16'sd373, 16'sd48, -16'sd607, -16'sd123, -16'sd1148, 16'sd383, 16'sd941, 16'sd213, -16'sd14},
'{-16'sd301, -16'sd754, -16'sd1979, 16'sd859, -16'sd1140, 16'sd583, -16'sd954, 16'sd679, -16'sd622, 16'sd425, -16'sd892, 16'sd84, 16'sd962, -16'sd331, 16'sd517, 16'sd680,16'sd252, -16'sd655, 16'sd1340, -16'sd683, -16'sd734, 16'sd1373, -16'sd723, -16'sd111, 16'sd119, 16'sd9, 16'sd250, -16'sd476, 16'sd26, 16'sd224, -16'sd36, -16'sd14,16'sd617, -16'sd810, -16'sd927, 16'sd504, -16'sd84, 16'sd298, -16'sd248, -16'sd19, 16'sd178, -16'sd441, -16'sd190, 16'sd502, 16'sd621, 16'sd985, -16'sd842, 16'sd562,16'sd458, 16'sd679, 16'sd279, -16'sd649, -16'sd1086, -16'sd201, 16'sd1127, 16'sd1253, -16'sd191, -16'sd925, 16'sd140, -16'sd498, 16'sd667, -16'sd309, -16'sd374, -16'sd636},
'{16'sd583, -16'sd456, 16'sd121, -16'sd600, 16'sd571, -16'sd439, 16'sd585, 16'sd182, 16'sd718, -16'sd477, -16'sd71, 16'sd133, 16'sd67, -16'sd1164, 16'sd295, -16'sd715,16'sd255, -16'sd237, 16'sd1385, 16'sd1760, -16'sd61, -16'sd866, 16'sd342, 16'sd763, 16'sd768, 16'sd1511, 16'sd357, -16'sd96, -16'sd1222, 16'sd719, -16'sd183, -16'sd190,16'sd360, -16'sd1396, -16'sd1356, 16'sd1204, 16'sd1341, 16'sd1685, -16'sd737, -16'sd29, -16'sd703, 16'sd165, 16'sd1276, 16'sd546, 16'sd1143, -16'sd965, -16'sd98, 16'sd563,16'sd176, 16'sd1409, -16'sd1039, -16'sd355, 16'sd780, 16'sd405, 16'sd339, -16'sd389, 16'sd475, -16'sd1324, -16'sd191, -16'sd392, -16'sd443, 16'sd1447, 16'sd669, -16'sd918},
'{16'sd480, -16'sd1087, -16'sd357, -16'sd844, -16'sd149, -16'sd165, 16'sd103, -16'sd201, 16'sd854, -16'sd1192, -16'sd669, 16'sd469, -16'sd742, 16'sd23, 16'sd477, 16'sd1006,16'sd245, 16'sd240, 16'sd1178, 16'sd1139, -16'sd324, 16'sd417, -16'sd816, 16'sd734, -16'sd336, -16'sd986, -16'sd349, 16'sd785, 16'sd670, 16'sd940, -16'sd1575, -16'sd916,16'sd416, -16'sd566, -16'sd869, 16'sd666, -16'sd438, -16'sd290, 16'sd587, -16'sd1644, -16'sd1359, -16'sd806, -16'sd1212, 16'sd632, 16'sd482, 16'sd955, -16'sd1678, 16'sd981,16'sd698, -16'sd594, -16'sd985, -16'sd329, 16'sd162, 16'sd1084, -16'sd667, 16'sd15, 16'sd764, 16'sd1174, -16'sd195, -16'sd649, 16'sd1090, 16'sd137, 16'sd397, 16'sd837},
'{16'sd670, -16'sd1081, -16'sd1074, 16'sd373, -16'sd893, -16'sd718, -16'sd1017, -16'sd318, -16'sd597, 16'sd876, -16'sd144, 16'sd960, -16'sd378, -16'sd429, 16'sd117, 16'sd737,16'sd18, -16'sd1036, -16'sd1501, -16'sd188, 16'sd627, -16'sd176, -16'sd1176, -16'sd104, -16'sd1674, -16'sd482, 16'sd1049, -16'sd117, 16'sd85, -16'sd170, -16'sd119, -16'sd160,16'sd2215, -16'sd469, -16'sd1014, 16'sd1703, 16'sd704, -16'sd134, -16'sd203, -16'sd509, 16'sd471, 16'sd336, 16'sd71, -16'sd61, 16'sd1026, -16'sd973, -16'sd604, -16'sd625,16'sd1405, -16'sd598, -16'sd82, 16'sd331, -16'sd781, -16'sd147, 16'sd1640, 16'sd558, 16'sd24, 16'sd288, 16'sd967, -16'sd1449, 16'sd939, -16'sd216, -16'sd819, 16'sd1434},
'{16'sd1166, -16'sd345, 16'sd421, -16'sd844, -16'sd446, 16'sd1474, 16'sd640, 16'sd970, -16'sd383, 16'sd662, 16'sd1155, -16'sd128, -16'sd528, -16'sd465, -16'sd158, 16'sd385,16'sd389, -16'sd424, 16'sd76, -16'sd1564, -16'sd137, -16'sd35, -16'sd625, 16'sd545, 16'sd23, 16'sd741, 16'sd818, 16'sd14, -16'sd482, -16'sd234, 16'sd513, 16'sd1777, -16'sd223,16'sd1109, -16'sd594, 16'sd72, -16'sd308, -16'sd1479, -16'sd43, 16'sd984, 16'sd664, -16'sd659, -16'sd933, 16'sd861, -16'sd495, 16'sd696, -16'sd184, 16'sd1069, 16'sd273,16'sd266, -16'sd547, -16'sd1261, -16'sd697, 16'sd878, 16'sd356, 16'sd1078, -16'sd808, -16'sd1069, 16'sd509, 16'sd668, -16'sd297, -16'sd1637, -16'sd591, -16'sd6},
'{-16'sd191, 16'sd867, 16'sd351, -16'sd89, -16'sd640, -16'sd136, 16'sd794, -16'sd6, -16'sd284, 16'sd42, -16'sd332, 16'sd616, 16'sd208, -16'sd582, 16'sd293, -16'sd1080,16'sd377, 16'sd1016, -16'sd1224, 16'sd9, -16'sd1181, -16'sd1204, 16'sd97, -16'sd904, 16'sd228, -16'sd24, 16'sd1256, 16'sd1069, 16'sd523, 16'sd1144, -16'sd523, -16'sd648,16'sd93, 16'sd701, 16'sd210, 16'sd81, -16'sd339, 16'sd123, 16'sd877, 16'sd569, 16'sd1028, -16'sd464, -16'sd197, -16'sd351, 16'sd72, -16'sd420, -16'sd968, -16'sd140,16'sd893, -16'sd748, 16'sd237, -16'sd145, -16'sd553, -16'sd59, 16'sd276, -16'sd13, 16'sd901, -16'sd392, -16'sd1801, -16'sd535, -16'sd195, -16'sd1386, 16'sd1006, 16'sd777},
'{16'sd626, 16'sd1427, -16'sd134, -16'sd163, -16'sd1199, 16'sd1192, 16'sd317, -16'sd801, -16'sd796, 16'sd196, -16'sd235, 16'sd18, 16'sd949, -16'sd363, -16'sd548, 16'sd1074,16'sd417, 16'sd270, -16'sd660, -16'sd246, -16'sd789, -16'sd993, -16'sd1024, -16'sd452, 16'sd1122, 16'sd563, 16'sd224, 16'sd3, 16'sd345, -16'sd1225, 16'sd374, -16'sd702,16'sd398, 16'sd484, 16'sd1412, -16'sd1271, 16'sd333, 16'sd299, -16'sd238, 16'sd53, 16'sd948, 16'sd639, -16'sd561, -16'sd1007, 16'sd664, -16'sd605, 16'sd0, 16'sd861,16'sd589, -16'sd11, 16'sd701, 16'sd186, 16'sd144, 16'sd470, 16'sd1383, 16'sd937, 16'sd25, -16'sd43, 16'sd531, -16'sd1375, -16'sd617, 16'sd2, 16'sd767, -16'sd880},
'{-16'sd731, 16'sd384, -16'sd1800, 16'sd695, 16'sd1837, -16'sd128, 16'sd1581, 16'sd725, -16'sd625, 16'sd556, 16'sd881, -16'sd222, 16'sd925, 16'sd375, -16'sd616, -16'sd1067,16'sd696, 16'sd7, -16'sd98, -16'sd1533, 16'sd147, 16'sd183, 16'sd1298, -16'sd530, -16'sd221, 16'sd169, 16'sd158, 16'sd257, -16'sd515, 16'sd246, -16'sd63, -16'sd395,16'sd263, -16'sd903, 16'sd67, -16'sd30, 16'sd938, -16'sd1321, -16'sd413, -16'sd630, 16'sd303, -16'sd61, -16'sd1220, -16'sd140, -16'sd223, 16'sd60, 16'sd1304, 16'sd1359,16'sd1004, -16'sd1669, 16'sd220, -16'sd69, -16'sd412, 16'sd347, 16'sd368, 16'sd1467, 16'sd310, -16'sd36, 16'sd723, 16'sd642, 16'sd753, 16'sd328, 16'sd1313, -16'sd473},
'{-16'sd1031, -16'sd684, 16'sd1000, 16'sd121, -16'sd489, 16'sd988, 16'sd1524, 16'sd374, -16'sd1356, -16'sd15, -16'sd369, -16'sd1454, -16'sd433, 16'sd193, 16'sd339, -16'sd1015,16'sd163, -16'sd242, 16'sd407, -16'sd781, -16'sd1876, -16'sd317, 16'sd198, 16'sd922, -16'sd67, 16'sd64, -16'sd85, 16'sd309, 16'sd324, -16'sd469, -16'sd341, 16'sd359,16'sd809, -16'sd915, -16'sd928, 16'sd914, -16'sd204, -16'sd1209, 16'sd750, 16'sd1, -16'sd310, -16'sd675, 16'sd175, 16'sd399, -16'sd389, -16'sd1498, 16'sd797, -16'sd516,16'sd16, -16'sd642, 16'sd255, -16'sd673, 16'sd1342, 16'sd979, 16'sd2067, 16'sd465, -16'sd320, 16'sd1170, 16'sd167, -16'sd569, 16'sd567, 16'sd685, -16'sd284, -16'sd96},
'{-16'sd166, -16'sd203, -16'sd492, 16'sd968, 16'sd292, 16'sd133, 16'sd385, 16'sd859, -16'sd924, -16'sd191, 16'sd179, -16'sd418, -16'sd836, 16'sd57, -16'sd929, 16'sd426,16'sd312, 16'sd1096, 16'sd7, -16'sd633, -16'sd730, 16'sd484, -16'sd525, 16'sd244, 16'sd577, -16'sd387, -16'sd537, 16'sd819, 16'sd531, -16'sd643, 16'sd2159, -16'sd281,16'sd204, -16'sd127, 16'sd718, -16'sd1026, -16'sd910, 16'sd523, 16'sd22, -16'sd1010, -16'sd338, -16'sd1332, 16'sd404, -16'sd728, -16'sd755, 16'sd1, -16'sd589, -16'sd13,16'sd71, 16'sd688, -16'sd573, 16'sd278, 16'sd83, -16'sd848, 16'sd295, 16'sd383, -16'sd651, 16'sd757, -16'sd484, -16'sd184, -16'sd339, 16'sd399, 16'sd1277, -16'sd603},
'{-16'sd1039, -16'sd756, -16'sd495, 16'sd726, -16'sd396, -16'sd530, -16'sd552, -16'sd203, -16'sd112, -16'sd1563, 16'sd926, -16'sd1511, 16'sd786, 16'sd91, -16'sd812, -16'sd1217,16'sd290, -16'sd589, -16'sd603, 16'sd706, 16'sd459, -16'sd115, -16'sd455, 16'sd427, 16'sd1097, 16'sd181, 16'sd229, 16'sd386, 16'sd314, 16'sd554, -16'sd196, 16'sd587, -16'sd486,16'sd1102, -16'sd176, 16'sd736, 16'sd1024, -16'sd337, 16'sd218, 16'sd627, -16'sd683, -16'sd367, -16'sd1567, -16'sd461, -16'sd631, -16'sd723, -16'sd261, -16'sd1127, -16'sd1396,16'sd402, 16'sd1013, -16'sd355, 16'sd466, 16'sd1099, 16'sd769, -16'sd261, 16'sd440, -16'sd888, -16'sd625, -16'sd558, 16'sd222, -16'sd1156, -16'sd609, 16'sd1},
'{16'sd464, 16'sd143, 16'sd768, 16'sd1270, 16'sd637, -16'sd197, -16'sd230, -16'sd213, 16'sd441, -16'sd316, -16'sd1093, 16'sd144, 16'sd931, -16'sd363, 16'sd1731, -16'sd1054,16'sd18, 16'sd1568, -16'sd1365, -16'sd1485, 16'sd343, -16'sd476, -16'sd1338, -16'sd164, 16'sd601, -16'sd1073, 16'sd1147, 16'sd287, -16'sd465, -16'sd480, -16'sd964, -16'sd531,16'sd1663, 16'sd1052, -16'sd752, -16'sd745, -16'sd410, -16'sd1209, 16'sd1490, -16'sd373, 16'sd548, -16'sd393, -16'sd102, -16'sd324, -16'sd637, -16'sd794, -16'sd162, -16'sd709,16'sd318, 16'sd972, -16'sd297, -16'sd778, 16'sd329, -16'sd334, -16'sd29, -16'sd397, 16'sd280, -16'sd237, 16'sd1138, -16'sd348, 16'sd510, -16'sd181, -16'sd631, 16'sd136},
'{16'sd357, -16'sd557, -16'sd79, 16'sd257, 16'sd752, 16'sd704, 16'sd434, 16'sd1020, -16'sd595, 16'sd122, -16'sd193, 16'sd181, 16'sd224, 16'sd777, 16'sd876, -16'sd214, 16'sd29, -16'sd953, -16'sd775, 16'sd142, -16'sd1097, -16'sd826, -16'sd478, -16'sd388, 16'sd200, 16'sd1045, 16'sd259, -16'sd136, 16'sd166, -16'sd13, -16'sd542, 16'sd630, 16'sd832, 16'sd380, 16'sd120, -16'sd219, -16'sd736, -16'sd74, 16'sd263, 16'sd140, -16'sd709, 16'sd1009, -16'sd351, -16'sd1336, -16'sd141, -16'sd563, -16'sd862, -16'sd404, -16'sd606, -16'sd752, 16'sd343, 16'sd708, -16'sd339, 16'sd534, 16'sd1054, -16'sd351, -16'sd470, -16'sd360, -16'sd560, 16'sd954, -16'sd1491, -16'sd277, -16'sd1309, -16'sd972},
'{16'sd234, -16'sd716, 16'sd674, -16'sd3, 16'sd299, -16'sd126, 16'sd1134, 16'sd950, -16'sd1228, -16'sd448, 16'sd276, -16'sd1061, 16'sd739, -16'sd876, 16'sd479, -16'sd1023, 16'sd1281, -16'sd1108, -16'sd405, 16'sd419, -16'sd158, 16'sd804, 16'sd660, -16'sd1329, 16'sd67, -16'sd565, 16'sd1437, 16'sd3, 16'sd780, 16'sd97, 16'sd575, -16'sd1410, 16'sd131, 16'sd632, -16'sd1172, 16'sd468, 16'sd780, 16'sd765, -16'sd1064, 16'sd191, -16'sd502, -16'sd1010, 16'sd363, -16'sd249, -16'sd747, -16'sd223, 16'sd159, 16'sd1248, 16'sd47, 16'sd394, -16'sd1424, -16'sd203, 16'sd853, -16'sd1534, 16'sd1073, 16'sd753, -16'sd162, -16'sd140, 16'sd426, 16'sd920, 16'sd1299, -16'sd740, -16'sd949, 16'sd1052},
'{16'sd559, 16'sd1534, -16'sd905, 16'sd989, -16'sd2311, -16'sd773, 16'sd1809, 16'sd799, 16'sd292, -16'sd622, 16'sd620, 16'sd77, -16'sd629, -16'sd508, -16'sd30, -16'sd344, -16'sd270, -16'sd81, -16'sd76, 16'sd267, -16'sd382, -16'sd215, -16'sd788, 16'sd569, -16'sd163, -16'sd1331, -16'sd88, 16'sd168, 16'sd886, 16'sd107, 16'sd205, 16'sd784, -16'sd96, 16'sd739, 16'sd623, 16'sd1033, 16'sd294, -16'sd1003, -16'sd549, -16'sd69, -16'sd377, -16'sd1169, 16'sd539, 16'sd209, 16'sd536, 16'sd48, -16'sd663, -16'sd201, 16'sd309, 16'sd313, 16'sd790, -16'sd813, 16'sd178, -16'sd140, 16'sd7, -16'sd1135, 16'sd406, -16'sd501, 16'sd582, -16'sd12, 16'sd438, -16'sd586, -16'sd171, -16'sd484},
'{-16'sd1263, 16'sd108, 16'sd1078, -16'sd6, 16'sd561, -16'sd804, 16'sd5, -16'sd1017, 16'sd289, 16'sd578, -16'sd484, -16'sd32, 16'sd274, 16'sd1310, -16'sd1023, -16'sd501, -16'sd10, 16'sd272, 16'sd917, -16'sd805, -16'sd1283, -16'sd360, -16'sd86, -16'sd1602, 16'sd215, -16'sd389, -16'sd261, -16'sd385, -16'sd1140, 16'sd665, -16'sd725, 16'sd315, 16'sd419, 16'sd563, 16'sd153, -16'sd691, -16'sd329, 16'sd441, 16'sd996, 16'sd125, -16'sd789, 16'sd464, 16'sd429, -16'sd606, 16'sd45, 16'sd710, 16'sd1899, 16'sd557, -16'sd1139, -16'sd127, 16'sd219, 16'sd127, -16'sd917, 16'sd984, -16'sd1219, 16'sd512, 16'sd1568, -16'sd423, -16'sd1066, 16'sd842, -16'sd174, -16'sd853, 16'sd2213, 16'sd510},
'{16'sd433, 16'sd96, 16'sd1385, -16'sd786, 16'sd147, -16'sd652, 16'sd322, 16'sd148, -16'sd1331, 16'sd291, -16'sd452, 16'sd275, 16'sd8, -16'sd369, -16'sd37, 16'sd236, 16'sd154, -16'sd756, -16'sd309, 16'sd425, -16'sd500, -16'sd233, 16'sd177, -16'sd1057, 16'sd89, 16'sd448, -16'sd216, 16'sd1024, 16'sd924, 16'sd1031, -16'sd832, 16'sd684, 16'sd1443, -16'sd1106, 16'sd532, 16'sd1136, -16'sd300, 16'sd671, -16'sd37, -16'sd758, 16'sd731, -16'sd227, -16'sd612, -16'sd519, -16'sd709, 16'sd1356, 16'sd251, 16'sd923, -16'sd30, -16'sd676, -16'sd618, -16'sd449, 16'sd819, 16'sd255, 16'sd709, -16'sd853, 16'sd1235, 16'sd123, 16'sd159, -16'sd860, 16'sd189, -16'sd168, -16'sd1139, -16'sd410},
'{-16'sd803, -16'sd468, -16'sd578, -16'sd1382, 16'sd137, -16'sd236, 16'sd1019, 16'sd472, -16'sd1275, 16'sd606, -16'sd247, 16'sd173, -16'sd429, -16'sd106, -16'sd314, -16'sd803, -16'sd1187, -16'sd355, 16'sd987, -16'sd287, 16'sd565, -16'sd1294, 16'sd108, -16'sd362, -16'sd1080, 16'sd123, 16'sd738, 16'sd693, 16'sd1323, -16'sd1976, -16'sd287, 16'sd564, 16'sd1076, -16'sd702, -16'sd821, -16'sd224, 16'sd840, -16'sd932, 16'sd550, -16'sd690, -16'sd3, 16'sd540, 16'sd47, -16'sd1796, 16'sd88, 16'sd195, -16'sd1328, 16'sd923, 16'sd476, 16'sd249, -16'sd360, -16'sd658, 16'sd397, 16'sd748, 16'sd335, 16'sd681, -16'sd703, -16'sd430, -16'sd616, 16'sd432, -16'sd414, -16'sd1648, 16'sd120, -16'sd137},
'{16'sd18, 16'sd905, 16'sd975, -16'sd206, 16'sd145, -16'sd1669, 16'sd937, -16'sd479, 16'sd1197, -16'sd448, 16'sd1155, 16'sd1322, -16'sd159, 16'sd742, -16'sd622, -16'sd154, -16'sd657, 16'sd267, 16'sd414, 16'sd861, -16'sd292, 16'sd119, 16'sd948, 16'sd37, -16'sd529, 16'sd106, 16'sd148, 16'sd863, -16'sd126, -16'sd807, -16'sd1949, 16'sd225, 16'sd65, -16'sd1127, -16'sd170, -16'sd109, 16'sd360, 16'sd220, 16'sd11, 16'sd713, -16'sd1300, -16'sd520, 16'sd721, 16'sd606, 16'sd533, -16'sd82, -16'sd874, 16'sd18, 16'sd920, -16'sd653, 16'sd388, -16'sd471, 16'sd35, 16'sd1013, 16'sd157, 16'sd93, -16'sd900, 16'sd125, -16'sd313, -16'sd1125, 16'sd564, 16'sd19, -16'sd486, -16'sd231},
'{16'sd135, 16'sd1134, 16'sd42, -16'sd6, 16'sd60, 16'sd819, -16'sd463, 16'sd1330, -16'sd541, 16'sd1541, -16'sd158, 16'sd1154, -16'sd230, -16'sd438, -16'sd1344, -16'sd414, -16'sd707, 16'sd497, 16'sd95, -16'sd665, 16'sd340, 16'sd265, 16'sd239, 16'sd446, -16'sd279, -16'sd596, -16'sd854, 16'sd1174, -16'sd648, 16'sd127, -16'sd149, 16'sd494, 16'sd658, 16'sd1007, -16'sd551, 16'sd921, 16'sd89, -16'sd286, -16'sd413, -16'sd342, 16'sd1274, 16'sd955, 16'sd946, -16'sd1171, -16'sd1075, -16'sd1128, 16'sd928, -16'sd38, -16'sd1784, -16'sd673, 16'sd532, -16'sd1102, 16'sd31, -16'sd260, 16'sd240, 16'sd1067, -16'sd2069, 16'sd1198, -16'sd291, 16'sd928, 16'sd528, -16'sd1735, 16'sd232, -16'sd15},
'{-16'sd1024, -16'sd69, 16'sd930, 16'sd498, 16'sd1349, 16'sd270, 16'sd1292, -16'sd92, 16'sd371, 16'sd667, 16'sd267, 16'sd928, 16'sd1324, -16'sd1543, -16'sd885, -16'sd676, -16'sd1172, -16'sd724, 16'sd56, 16'sd502, -16'sd1425, -16'sd931, 16'sd567, 16'sd567, 16'sd567, -16'sd318, 16'sd116, -16'sd1440, 16'sd1712, -16'sd823, 16'sd196, -16'sd888, -16'sd1304, 16'sd708, 16'sd143, 16'sd838, -16'sd1445, 16'sd439, 16'sd599, -16'sd1567, -16'sd878, -16'sd842, -16'sd226, 16'sd90, 16'sd243, -16'sd288, -16'sd1072, 16'sd1333, -16'sd254, 16'sd355, 16'sd958, 16'sd834, -16'sd285, -16'sd407, -16'sd1094, 16'sd1046, -16'sd343, 16'sd69, -16'sd164, 16'sd863, 16'sd1206, -16'sd960, 16'sd14, 16'sd171},
'{16'sd704, -16'sd363, -16'sd258, 16'sd1151, 16'sd346, -16'sd688, 16'sd176, -16'sd809, -16'sd1461, 16'sd1350, -16'sd1085, 16'sd1427, 16'sd871, -16'sd198, -16'sd33, -16'sd771, 16'sd332, 16'sd580, 16'sd1048, -16'sd1554, 16'sd653, 16'sd712, -16'sd844, 16'sd31, -16'sd791, -16'sd442, 16'sd1139, -16'sd3, 16'sd735, -16'sd405, 16'sd75, -16'sd674, -16'sd337, -16'sd440, 16'sd262, -16'sd274, -16'sd364, -16'sd1573, 16'sd919, -16'sd1525, 16'sd271, 16'sd214, 16'sd162, -16'sd537, 16'sd253, 16'sd351, 16'sd1081, -16'sd214, 16'sd440, -16'sd261, -16'sd493, -16'sd1191, 16'sd286, -16'sd167, -16'sd44, 16'sd131, -16'sd115, 16'sd1476, -16'sd436, 16'sd613, 16'sd296, 16'sd1009, -16'sd875, -16'sd1197},
'{16'sd50, 16'sd904, 16'sd233, -16'sd32, 16'sd975, -16'sd679, -16'sd1149, 16'sd1388, -16'sd1231, 16'sd305, 16'sd441, 16'sd41, -16'sd128, -16'sd390, 16'sd987, 16'sd971, 16'sd574, 16'sd1098, 16'sd403, -16'sd301, -16'sd82, -16'sd591, 16'sd522, 16'sd49, -16'sd1132, -16'sd526, 16'sd1289, -16'sd274, -16'sd143, 16'sd439, -16'sd1385, 16'sd765, -16'sd486, 16'sd755, -16'sd175, 16'sd333, 16'sd1168, 16'sd35, 16'sd640, 16'sd1749, 16'sd252, 16'sd1119, -16'sd1198, 16'sd132, -16'sd82, -16'sd563, -16'sd1891, 16'sd309, -16'sd1099, -16'sd139, 16'sd106, -16'sd46, 16'sd48, 16'sd745, 16'sd392, -16'sd623, -16'sd1252, 16'sd139, 16'sd474, -16'sd201, 16'sd689, 16'sd453, 16'sd212, -16'sd179},
'{16'sd293, -16'sd111, 16'sd173, -16'sd150, 16'sd270, 16'sd1211, -16'sd443, -16'sd1279, 16'sd1193, 16'sd264, 16'sd5, -16'sd1593, -16'sd357, -16'sd1274, -16'sd1445, 16'sd407, -16'sd136, -16'sd753, 16'sd758, 16'sd603, -16'sd521, -16'sd597, -16'sd1103, -16'sd1285, -16'sd502, 16'sd469, 16'sd151, -16'sd1057, -16'sd796, 16'sd698, -16'sd512, 16'sd1782, -16'sd673, -16'sd337, -16'sd1676, -16'sd376, -16'sd216, 16'sd1264, -16'sd359, 16'sd359, -16'sd481, 16'sd625, -16'sd6, -16'sd152, -16'sd534, 16'sd1641, -16'sd721, 16'sd171, -16'sd106, 16'sd867, 16'sd451, -16'sd70, -16'sd469, 16'sd1933, 16'sd398, -16'sd520, -16'sd712, -16'sd38, -16'sd1149, -16'sd569, -16'sd980, 16'sd449, 16'sd421, -16'sd1001},
'{-16'sd883, -16'sd722, 16'sd831, 16'sd306, 16'sd991, -16'sd996, 16'sd670, 16'sd456, 16'sd222, 16'sd455, -16'sd648, -16'sd53, -16'sd368, 16'sd214, -16'sd810, -16'sd654, 16'sd773, 16'sd491, -16'sd568, -16'sd122, 16'sd631, 16'sd227, 16'sd502, 16'sd1156, -16'sd473, 16'sd541, -16'sd313, 16'sd684, 16'sd160, -16'sd4, 16'sd469, -16'sd196, 16'sd1032, -16'sd791, -16'sd213, 16'sd520, 16'sd779, 16'sd439, -16'sd478, -16'sd702, 16'sd168, 16'sd75, 16'sd468, 16'sd1154, 16'sd1442, -16'sd463, -16'sd92, 16'sd221, 16'sd144, -16'sd308, 16'sd1026, 16'sd654, -16'sd56, -16'sd1493, -16'sd177, -16'sd2581, 16'sd1084, 16'sd252, 16'sd296, 16'sd1312, 16'sd367, 16'sd270, -16'sd294, -16'sd920},
'{-16'sd1286, -16'sd863, -16'sd934, 16'sd73, 16'sd76, 16'sd565, -16'sd66, 16'sd770, -16'sd42, 16'sd190, -16'sd650, 16'sd206, -16'sd503, -16'sd964, -16'sd631, -16'sd453, -16'sd1410, -16'sd606, -16'sd715, -16'sd674, 16'sd304, -16'sd1468, 16'sd827, -16'sd554, -16'sd731, -16'sd1044, -16'sd837, -16'sd323, 16'sd138, -16'sd1036, 16'sd1167, 16'sd555, -16'sd17, -16'sd865, -16'sd1062, -16'sd231, 16'sd1195, -16'sd592, 16'sd675, -16'sd993, -16'sd638, -16'sd169, -16'sd556, 16'sd841, -16'sd869, 16'sd378, 16'sd897, 16'sd507, -16'sd475, 16'sd160, 16'sd141, -16'sd74, -16'sd887, -16'sd13, 16'sd690, 16'sd368, 16'sd34, -16'sd833, 16'sd1350, -16'sd1018, -16'sd368, 16'sd2, 16'sd744, 16'sd975},
'{16'sd526, -16'sd727, 16'sd688, 16'sd300, -16'sd239, -16'sd991, 16'sd958, -16'sd1463, 16'sd564, -16'sd511, 16'sd298, 16'sd118, -16'sd664, 16'sd840, 16'sd1010, -16'sd855, 16'sd120, 16'sd306, -16'sd1049, -16'sd1045, -16'sd89, 16'sd565, 16'sd600, -16'sd373, 16'sd35, 16'sd642, 16'sd518, -16'sd39, 16'sd328, -16'sd284, 16'sd10, 16'sd713, -16'sd619, 16'sd1133, -16'sd923, -16'sd742, 16'sd798, -16'sd975, -16'sd737, 16'sd513, -16'sd29, 16'sd584, 16'sd2121, 16'sd305, -16'sd12, -16'sd497, 16'sd132, -16'sd1029, 16'sd1182, -16'sd262, 16'sd53, -16'sd953, -16'sd130, -16'sd608, 16'sd352, 16'sd561, -16'sd8, -16'sd166, -16'sd1289, -16'sd332, 16'sd443, 16'sd1143, -16'sd733, -16'sd738},
'{16'sd598, -16'sd405, 16'sd519, 16'sd1306, 16'sd427, 16'sd1274, 16'sd195, -16'sd709, -16'sd312, -16'sd1807, 16'sd696, 16'sd289, -16'sd139, 16'sd1096, -16'sd1021, -16'sd791, 16'sd1334, 16'sd6, 16'sd1195, -16'sd1060, -16'sd870, -16'sd582, -16'sd195, 16'sd638, -16'sd785, 16'sd872, -16'sd60, -16'sd283, -16'sd338, -16'sd405, 16'sd211, -16'sd366, -16'sd803, 16'sd765, -16'sd530, 16'sd1186, -16'sd349, 16'sd890, 16'sd265, -16'sd128, -16'sd401, 16'sd934, -16'sd1009, 16'sd192, 16'sd68, -16'sd295, -16'sd436, -16'sd211, 16'sd974, -16'sd345, 16'sd811, 16'sd1336, 16'sd7, 16'sd158, -16'sd994, 16'sd887, -16'sd1239, 16'sd224, 16'sd1444, 16'sd987, 16'sd997, -16'sd313, -16'sd297, -16'sd893  }

};


typedef logic signed [15:0] signed_matrix_1x32_t[32];

const signed_matrix_1x32_t biases_2 = '{-16'sd1, -16'sd6, -16'sd4, 16'sd4, -16'sd6, 16'sd8, -16'sd2, -16'sd1, -16'sd3, 16'sd4, 16'sd3, -16'sd4, -16'sd3, 16'sd8, -16'sd3, -16'sd1, -16'sd6, -16'sd6, 16'sd0, 16'sd5, 16'sd2, -16'sd2, 16'sd0, 16'sd3, -16'sd3, 16'sd1, 16'sd2, 16'sd3, 16'sd14, -16'sd2, 16'sd1, 16'sd4};

integer i, j;
logic signed [31:0] sum; // 用于累加，扩展位宽以避免溢出


logic signed [15:0] temp_output_data[0:31]; // 临时存储调整后的结果

always @(posedge clk or posedge reset) begin
    if (reset) begin
        for (i = 0; i < 32; i = i + 1) begin
            output_data[i] <= 0; // 在复位时清零输出数据
        end
        valid_out <= 0; // 重置时，输出数据无效
    end else if (valid_in) begin
        for (i = 0; i < 32; i = i + 1) begin
            sum = 0; // 在开始累加前初始化sum为0
            for (j = 0; j < 64; j = j + 1) begin
                // 执行矩阵乘法和累加
                sum = sum + (input_data[j] * weights_2[i][j]);
            end
            // 所有加权和完成后，整体右移12位来调整格式
            sum = sum >>> 12;
            sum = sum + biases_2[i]; // 加上偏置
            temp_output_data[i] = sum[15:0]; // 临时存储调整后的结果
        end
        // 使用单独的循环将临时结果赋值给输出，确保使用非阻塞性赋值
        for (i = 0; i < 32; i = i + 1) begin
            output_data[i] <= temp_output_data[i];
        end
        valid_out <= 1; // 处理完成后，标记输出数据为有效
    end
end


assign ready_out = 1;



endmodule